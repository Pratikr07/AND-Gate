`timescale 1ns/1ns
module tb_and_gate;

   reg a,b;
   wire y;

   and_gate uut(.a(a),.b(b),.y(y));

   initial 
   begin
      $dumpfile("and.vcd");
      $dumpvars(0,tb_and_gate);

      a=0; b=0; #10;
      a=0; b=1; #10;
      a=1; b=0; #10;
      a=1; b=1; #10;

      $finish;
   end
endmodule
